library IEEE;
use IEEE.std_logic_1164.all; 
use IEEE.numeric_std.all; 
use types.all;

entity CONNECTED is
	generic(
		INSTRUCTION_SIZE: INTEGER := 16
	);						   
	port(	 													
		RESET: in STD_LOGIC;
		CLK: in STD_LOGIC;	
		
		REG_MATRIX: out matrix8(15 downto 0)
	);

end entity CONNECTED;

architecture CONNECTED_ARCHITECTURE of CONNECTED is

--
-- Component declaration
--

component REGISTERS_BLACK_BOX is
	generic(
		NR_BITS: INTEGER:= 8;
		NR_OF_REGISTERS: INTEGER:= 16
	);
	port(	   
		RESET: in STD_LOGIC;
		ENABLE: in STD_LOGIC;
		CLK: in STD_LOGIC;
		
		REGISTER_UPDATE_INPUT: in STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);
		
		FIRST_MUX_SEL: in INTEGER;
		SECOND_MUX_SEL: in INTEGER;
		
		FIRST_REGISTER_OUT: out STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);
		SECOND_REGISTER_OUT: out STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);
		
		REGISTER_MATRIX_OUT: out matrix8(15 downto 0)
	);
end component REGISTERS_BLACK_BOX;

component ALU_BLACK_BOX is										  
	generic(
		NR_BITS: INTEGER := 8;
		INPUT_MUX_SEL_NUMBER: INTEGER := 2;
		OUTPUT_MUX_SEL_NUMBER: INTEGER := 18
	);
	port( 
		FIRST_REGISTER_INPUT: in STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);
		SECOND_REGISTER_INPUT: in STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);
		CONSTANT_INPUT: in STD_LOGIC_VECTOR(NR_BITS - 1 downto 0); 
		
		SEL_MUX_INPUT: in INTEGER;	 	--muxul care alege registru/constanta
		SEL_MUX_OUTPUT: in INTEGER;	    --muxul care alege operatia care iese
		
		ZERO_FLAG: inout STD_LOGIC;
		CARRY_FLAG: inout STD_LOGIC;
		
		RESULT_OUTPUT: out STD_LOGIC_VECTOR(NR_BITS - 1 downto 0)
	);
end component ALU_BLACK_BOX; 

component DECODER_BLACK_BOX is
	generic(
		NR_BITS: INTEGER := 8; 			 
		INSTRUCTION_BITS: INTEGER := 16
	);						   
	port(
		INSTRUCTION: in STD_LOGIC_VECTOR(INSTRUCTION_BITS - 1 downto 0);
		
		CONSTANT_NUMBER: out STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);
		REGISTER_FIRST_NUMBER: out INTEGER;	
		REGISTER_SECOND_NUMBER: out INTEGER;
		
		REG_ENABLE: out STD_LOGIC;				--0 - daca e jump/call etc 
		
		ALU_INPUT_SEL: out INTEGER;
		ALU_OUTPUT_SEL: out INTEGER;
		
		FLOW_MODE: out INTEGER;
		FLOW_LOAD: out INTEGER;
		
		FLOW_COND: out INTEGER;
		FLOW_SEL: out INTEGER;	
		
		ZERO_FLAG: in STD_LOGIC;
		CARRY_FLAG: in STD_LOGIC
	);								
end component DECODER_BLACK_BOX;

component COUNTER_BLACK_BOX is		
	generic(
		MODULO: INTEGER := 254
	);
	port(
		CLK: in STD_LOGIC;	 
		MODE: in INTEGER;	--0 numara, 1 load
		PARALLEL_LOAD: in INTEGER;
		RESET: in STD_LOGIC;
	    OUTPUT: inout INTEGER
	);
end component COUNTER_BLACK_BOX;

component ROM is
	generic(
		NR_ADDRESSES:INTEGER := 256;
		WORD_LEN: INTEGER:= 16
	);						   
	port(
		ADDRESS: in INTEGER;
		OUTPUT: out STD_LOGIC_VECTOR(WORD_LEN - 1 downto 0)
	);
end component ROM;

component CLK_DIVIDER is
	port(
		CLK: in STD_LOGIC;
		CLK_REGISTER: out STD_LOGIC;
		CLK_COUNTER: out STD_LOGIC
	);
end component CLK_DIVIDER;	  

component FLOW_BLACK_BOX is  
	port(	  				
		MODE: in INTEGER;
		LOAD: in INTEGER; 
		
		COND: in INTEGER;
		SEL: in INTEGER;
		
		ZERO: in STD_LOGIC;
		CARRY: in STD_LOGIC;
		
		MODE_OUT: out INTEGER;
		LOAD_OUT: out INTEGER
	);
end component FLOW_BLACK_BOX;							   						   		

--
-- Signal declaration
--

signal FLOW_MODE: INTEGER := 0;
signal FLOW_LOAD: INTEGER := 0;

--signal COUNTER_MODE: INTEGER := 0;
--signal COUNTER_PARALLEL_LOAD: INTEGER := 0;	
signal COUNTER_OUTPUT: INTEGER;

signal CLK_REGISTER: STD_LOGIC;
signal CLK_COUNTER: STD_LOGIC;

signal ROM_INSTRUCTION: STD_LOGIC_VECTOR(15 downto 0);

signal DECODER_CONSTANT_NUMBER: STD_LOGIC_VECTOR(7 downto 0);
signal DECODER_REGISTER_FIRST_NUMBER: INTEGER;
signal DECODER_REGISTER_SECOND_NUMBER: INTEGER;
signal DECODER_REG_ENABLE: STD_LOGIC := '1';
signal DECODER_ALU_INPUT_SEL: INTEGER;
signal DECODER_ALU_OUTPUT_SEL: INTEGER;	
signal DECODER_FLOW_MODE: INTEGER;
signal DECODER_FLOW_LOAD: INTEGER; 
signal DECODER_FLOW_COND: INTEGER;
signal DECODER_FLOW_SEL: INTEGER;

signal REGISTER_FIRST_REGISTER_OUT: STD_LOGIC_VECTOR(7 downto 0);
signal REGISTER_SECOND_REGISTER_OUT: STD_LOGIC_VECTOR(7 downto 0);


signal FLAGS_ZERO_FLAG: STD_LOGIC := '0';
signal FLAGS_CARRY_FLAG: STD_LOGIC := '0';

signal ALU_RESULT_OUTPUT: STD_LOGIC_VECTOR(7 downto 0);	 

begin
	ALU_TAG: ALU_BLACK_BOX port map(
		REGISTER_FIRST_REGISTER_OUT,
		REGISTER_SECOND_REGISTER_OUT,
		DECODER_CONSTANT_NUMBER,
		DECODER_ALU_INPUT_SEL,
		DECODER_ALU_OUTPUT_SEL,
		FLAGS_ZERO_FLAG,
		FLAGS_CARRY_FLAG,
		ALU_RESULT_OUTPUT
	);
	DECODER_TAG: DECODER_BLACK_BOX port map(
		ROM_INSTRUCTION,
		DECODER_CONSTANT_NUMBER,
		DECODER_REGISTER_FIRST_NUMBER,
		DECODER_REGISTER_SECOND_NUMBER,
		DECODER_REG_ENABLE,
		DECODER_ALU_INPUT_SEL,
		DECODER_ALU_OUTPUT_SEL,
		DECODER_FLOW_MODE,
		DECODER_FLOW_LOAD,
		DECODER_FLOW_COND,
		DECODER_FLOW_SEL,
		FLAGS_ZERO_FLAG,
		FLAGS_CARRY_FLAG
	);					  
	REGISTER_TAG: REGISTERS_BLACK_BOX port map(
		RESET,
		DECODER_REG_ENABLE,
		CLK_REGISTER,
		ALU_RESULT_OUTPUT,
		DECODER_REGISTER_FIRST_NUMBER,
		DECODER_REGISTER_SECOND_NUMBER,
		REGISTER_FIRST_REGISTER_OUT,
		REGISTER_SECOND_REGISTER_OUT,
		REG_MATRIX
	);	
	CLK_DIVIDER_TAG: CLK_DIVIDER port map(
		CLK,
		CLK_REGISTER,
		CLK_COUNTER
	);
	COUNTER_TAG: COUNTER_BLACK_BOX port map(
		CLK_COUNTER,
		FLOW_MODE,
		FLOW_LOAD,
		RESET,
		COUNTER_OUTPUT
	);
	ROM_TAG: ROM port map(
		COUNTER_OUTPUT,
		ROM_INSTRUCTION
	);	
	FLOW_TAG: FLOW_BLACK_BOX port map( 
		DECODER_FLOW_MODE,
		DECODER_FLOW_LOAD, 
		DECODER_FLOW_COND,
		DECODER_FLOW_SEL,
		FLAGS_ZERO_FLAG,
		FLAGS_CARRY_FLAG,
		FLOW_MODE,
		FLOW_LOAD
	);	 
end architecture CONNECTED_ARCHITECTURE;