library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use types.all;

entity ALU_BLACK_BOX is										  
	generic(
		NR_BITS: INTEGER := 8;
		INPUT_MUX_SEL_NUMBER: INTEGER := 2;
		OUTPUT_MUX_SEL_NUMBER: INTEGER := 18
	);
	port( 
		FIRST_REGISTER_INPUT: in STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);
		SECOND_REGISTER_INPUT: in STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);
		CONSTANT_INPUT: in STD_LOGIC_VECTOR(NR_BITS - 1 downto 0); 
		
		SEL_MUX_INPUT: in INTEGER;	 	--muxul care alege registru/constanta
		SEL_MUX_OUTPUT: in INTEGER;	    --muxul care alege operatia care iese
		
		ZERO_FLAG: inout STD_LOGIC;
		CARRY_FLAG: inout STD_LOGIC;
		
		RESULT_OUTPUT: out STD_LOGIC_VECTOR(NR_BITS - 1 downto 0)
	);
end entity ALU_BLACK_BOX;									  

architecture ALU_BLACK_BOX_ARCHITECTURE of ALU_BLACK_BOX is

component MUX_INPUT is 	
	generic(
		NR_INPUTS: INTEGER := 2;	--0 - registru; 1 - constanta						 
		NR_BITS: INTEGER := 8
		);
	port(
		INPUT_MATRIX: in matrix(NR_INPUTS - 1 downto 0);
		SELECTION: in INTEGER;
		OUTPUT: out STD_LOGIC_VECTOR(NR_BITS - 1 downto 0)
	);
end component;


component ADD is
	generic(
		NR_BITS: INTEGER := 8
	);
	port(
		FIRST_NUMBER:in STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);
		SECOND_NUMBER:in STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);
		RESULT:out STD_LOGIC_VECTOR(NR_BITS - 1 downto 0); 
		ZERO_FLAG: out STD_LOGIC;
		CARRY:out STD_LOGIC
	);
end component; 

component ADDCY is
	generic(
		NR_BITS: INTEGER := 8
	);
	port(
		FIRST_NUMBER: in STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);
		SECOND_NUMBER: in STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);
		CARRY_IN: in STD_LOGIC;
		CARRY_OUT: out STD_LOGIC;	
		ZERO_FLAG: out STD_LOGIC;
		RESULT: out STD_LOGIC_VECTOR(NR_BITS - 1 downto 0)
	);
end component;

component ANDD is
	generic(
		NR_BITS: INTEGER := 8
	);						  
	port(
	FIRST_NUMBER: in STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);
	SECOND_NUMBER: in STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);
	RESULT: inout STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);
	ZERO_FLAG: out STD_LOGIC
	);
end component;	

component ORR is
	generic(
		NR_BITS: INTEGER := 8
	);						 
	port(
		FIRST_NUMBER: in STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);
		SECOND_NUMBER: in STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);
		RESULT: out STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);
		ZERO_FLAG: out STD_LOGIC
	);
end component;	

component SUB is
	generic(
		NR_BITS: INTEGER:= 8
	);							
	port(
		FIRST_NUMBER:in STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);
		SECOND_NUMBER: in STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);
		RESULT: out STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);	   
		ZERO_FLAG: out STD_LOGIC;
		BORROW: out STD_LOGIC
	);						
end component;	 

component SUBCY is
	generic(
		NR_BITS: INTEGER := 8
	);						  
	port(
		FIRST_NUMBER: in STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);
		SECOND_NUMBER: in STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);
		BORROW_IN: in STD_LOGIC;
		BORROW_OUT: out STD_LOGIC;						  
		ZERO_FLAG: out STD_LOGIC;
		RESULT: out STD_LOGIC_VECTOR(NR_BITS - 1 downto 0)
	);
end component;	

component XORR is
	generic(
		NR_BITS: INTEGER := 8
	);						 
	port(
		FIRST_NUMBER: in STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);
		SECOND_NUMBER: in STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);
		RESULT: out STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);
		ZERO_FLAG: out STD_LOGIC
	);
end component;

component SR0 is
	generic(
		NR_BITS:INTEGER := 8
	);						 
	port(
		FIRST_NUMBER:in STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);
		RESULT:out STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);	
		ZERO_FLAG: out STD_LOGIC;
		CARRY_FLAG: out STD_LOGIC
	);
end component;		

component SR1 is
	generic(
		NR_BITS:INTEGER := 8
	);						 
	port(
		FIRST_NUMBER:in STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);
		RESULT:out STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);	
		ZERO_FLAG: out STD_LOGIC;
		CARRY_FLAG: out STD_LOGIC
	);
end component SR1;	

component SRX is
	generic(
		NR_BITS:INTEGER := 8
	);						 
	port(
		FIRST_NUMBER:in STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);
		RESULT:out STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);	
		ZERO_FLAG: out STD_LOGIC;
		CARRY_FLAG: out STD_LOGIC
	);
end component SRX;	

component SRAA is
	generic(
		NR_BITS:INTEGER := 8
	);						 
	port(
		FIRST_NUMBER:in STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);
		CARRY_IN: in STD_LOGIC;
		RESULT:out STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);	
		ZERO_FLAG: out STD_LOGIC;
		CARRY_OUT: out STD_LOGIC
	);
end component SRAA;

component RR is
	generic(
		NR_BITS:INTEGER := 8
	);						 
	port(
		FIRST_NUMBER:in STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);
		RESULT:out STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);	
		ZERO_FLAG: out STD_LOGIC;
		CARRY_FLAG: out STD_LOGIC
	);
end component RR;		 

component SL0 is
	generic(
		NR_BITS:INTEGER := 8
	);						 
	port(
		FIRST_NUMBER:in STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);
		RESULT:out STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);	
		ZERO_FLAG: out STD_LOGIC;
		CARRY_FLAG: out STD_LOGIC
	);
end component SL0;		

component SL1 is
	generic(
		NR_BITS:INTEGER := 8
	);						 
	port(
		FIRST_NUMBER:in STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);
		RESULT:out STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);	
		ZERO_FLAG: out STD_LOGIC;
		CARRY_FLAG: out STD_LOGIC
	);
end component SL1;	 

component SLX is
	generic(
		NR_BITS:INTEGER := 8
	);						 
	port(
		FIRST_NUMBER:in STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);
		RESULT:out STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);	
		ZERO_FLAG: out STD_LOGIC;
		CARRY_FLAG: out STD_LOGIC
	);
end component SLX;		

component SLAA is
	generic(
		NR_BITS:INTEGER := 8
	);						 
	port(
		FIRST_NUMBER:in STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);
		CARRY_IN: in STD_LOGIC;
		RESULT:out STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);	
		ZERO_FLAG: out STD_LOGIC;
		CARRY_OUT: out STD_LOGIC
	);
end component SLAA;

component RL is
	generic(
		NR_BITS:INTEGER := 8
	);						 
	port(
		FIRST_NUMBER:in STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);
		RESULT:out STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);	
		ZERO_FLAG: out STD_LOGIC;
		CARRY_FLAG: out STD_LOGIC
	);
end component;	

component LOAD is 
	generic(
		NR_BITS: INTEGER := 8
	);						  
	port(
		FIRST_NUMBER: in STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);
		RESULT: out STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);
		ZERO_FLAG: out STD_LOGIC
	);
	
end component LOAD;

component MUX_OUTPUT is
	generic(
		NR_INPUTS: INTEGER := 18;	--18 operatii						 
		NR_BITS: INTEGER := 8
		);
		
	port(
		INPUT_MATRIX: in matrix(NR_INPUTS - 1 downto 0);
		SELECTION: in INTEGER;
		OUTPUT: out STD_LOGIC_VECTOR(NR_BITS - 1 downto 0)
	);
end component MUX_OUTPUT;

signal SECOND_OPERAND: STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);
signal AUXILIAR_MATRIX_INPUT: matrix(INPUT_MUX_SEL_NUMBER - 1 downto 0);	

signal ADD_RESULT:    STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);
signal ADDCY_RESULT:  STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);
signal AND_RESULT:    STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);
signal OR_RESULT:     STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);
signal SUB_RESULT:    STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);
signal SUBCY_RESULT:  STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);
signal XOR_RESULT:    STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);
signal SR0_RESULT:    STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);
signal SR1_RESULT:    STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);
signal SRX_RESULT:    STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);
signal SRA_RESULT:    STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);
signal RR_RESULT:     STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);
signal SL0_RESULT:    STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);
signal SL1_RESULT:    STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);
signal SLX_RESULT:    STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);
signal SLA_RESULT:    STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);
signal RL_RESULT:     STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);	  
signal LOAD_RESULT:   STD_LOGIC_VECTOR(NR_BITS - 1 downto 0);

signal ZERO_MATRIX:   STD_LOGIC_VECTOR(OUTPUT_MUX_SEL_NUMBER - 1 downto 0) := "000000000000000000";
signal CARRY_MATRIX:  STD_LOGIC_VECTOR(OUTPUT_MUX_SEL_NUMBER - 1 downto 0) := "000000000000000000";

signal AUXILIAR_MATRIX_OUTPUT: matrix(OUTPUT_MUX_SEL_NUMBER - 1 downto 0);

begin			
	AUXILIAR_MATRIX_INPUT(0) <= SECOND_REGISTER_INPUT;
	AUXILIAR_MATRIX_INPUT(1) <= CONSTANT_INPUT;
	FIRST_MUX_TAG: MUX_INPUT port map(AUXILIAR_MATRIX_INPUT, SEL_MUX_INPUT, SECOND_OPERAND);
	
	ADD_TAG:    ADD   port map(FIRST_REGISTER_INPUT, SECOND_OPERAND, ADD_RESULT, ZERO_MATRIX(0), CARRY_MATRIX(0));
	ADDCY_TAG:  ADDCY port map(FIRST_REGISTER_INPUT, SECOND_OPERAND, CARRY_MATRIX(1), CARRY_MATRIX(1), ZERO_MATRIX(1), ADDCY_RESULT);
	AND_TAG:    ANDD  port map(FIRST_REGISTER_INPUT, SECOND_OPERAND, AND_RESULT, ZERO_MATRIX(2));
	OR_TAG:     ORR   port map(FIRST_REGISTER_INPUT, SECOND_OPERAND, OR_RESULT, ZERO_MATRIX(3));
	SUB_TAG:    SUB   port map(FIRST_REGISTER_INPUT, SECOND_OPERAND, SUB_RESULT, ZERO_MATRIX(4), CARRY_MATRIX(4));
	SUBCY_TAG:  SUBCY port map(FIRST_REGISTER_INPUT, SECOND_OPERAND, CARRY_MATRIX(5), CARRY_MATRIX(5), ZERO_MATRIX(5), SUBCY_RESULT);
	XOR_TAG:    XORR  port map(FIRST_REGISTER_INPUT, SECOND_OPERAND, XOR_RESULT, ZERO_MATRIX(6));
	SR0_TAG:    SR0   port map(FIRST_REGISTER_INPUT, SR0_RESULT, ZERO_MATRIX(7), CARRY_MATRIX(7));
	SR1_TAG:    SR1   port map(FIRST_REGISTER_INPUT, SR1_RESULT, ZERO_MATRIX(8), CARRY_MATRIX(8));
	SRX_TAG:    SRX   port map(FIRST_REGISTER_INPUT, SRX_RESULT, ZERO_MATRIX(9), CARRY_MATRIX(9));
	SRA_TAG:    SRAA  port map(FIRST_REGISTER_INPUT, CARRY_MATRIX(10), SRA_RESULT, ZERO_MATRIX(10), CARRY_MATRIX(10));
	RR_TAG:     RR    port map(FIRST_REGISTER_INPUT, RR_RESULT, ZERO_MATRIX(11), CARRY_MATRIX(11));
	SL0_TAG:    SL0   port map(FIRST_REGISTER_INPUT, SL0_RESULT, ZERO_MATRIX(12), CARRY_MATRIX(12));
	SL1_TAG:    SL1   port map(FIRST_REGISTER_INPUT, SL1_RESULT, ZERO_MATRIX(13), CARRY_MATRIX(13));
	SLX_TAG:    SLX   port map(FIRST_REGISTER_INPUT, SLX_RESULT, ZERO_MATRIX(14), CARRY_MATRIX(14));
	SLA_TAG:    SLAA  port map(FIRST_REGISTER_INPUT, CARRY_FLAG, SLA_RESULT, ZERO_MATRIX(15), CARRY_MATRIX(15));
	RL_TAG:     RL    port map(FIRST_REGISTER_INPUT, RL_RESULT, ZERO_MATRIX(16), CARRY_MATRIX(16)); 
	LOAD_TAG:   LOAD  port map(SECOND_OPERAND, LOAD_RESULT, ZERO_MATRIX(17));
	
	AUXILIAR_MATRIX_OUTPUT(0)  <= ADD_RESULT;
	AUXILIAR_MATRIX_OUTPUT(1)  <= ADDCY_RESULT;	  
	AUXILIAR_MATRIX_OUTPUT(2)  <= AND_RESULT;
	AUXILIAR_MATRIX_OUTPUT(3)  <= OR_RESULT;
	AUXILIAR_MATRIX_OUTPUT(4)  <= SUB_RESULT;
	AUXILIAR_MATRIX_OUTPUT(5)  <= SUBCY_RESULT;
	AUXILIAR_MATRIX_OUTPUT(6)  <= XOR_RESULT;	  
	AUXILIAR_MATRIX_OUTPUT(7)  <= SR0_RESULT;
	AUXILIAR_MATRIX_OUTPUT(8)  <= SR1_RESULT;
	AUXILIAR_MATRIX_OUTPUT(9)  <= SRX_RESULT;
	AUXILIAR_MATRIX_OUTPUT(10) <= SRA_RESULT;
	AUXILIAR_MATRIX_OUTPUT(11) <= RR_RESULT;	  
	AUXILIAR_MATRIX_OUTPUT(12) <= SL0_RESULT;
	AUXILIAR_MATRIX_OUTPUT(13) <= SL1_RESULT;
	AUXILIAR_MATRIX_OUTPUT(14) <= SLX_RESULT;
	AUXILIAR_MATRIX_OUTPUT(15) <= SLA_RESULT;
	AUXILIAR_MATRIX_OUTPUT(16) <= RL_RESULT;
	AUXILIAR_MATRIX_OUTPUT(17) <= LOAD_RESULT;
	
	process(ZERO_MATRIX, CARRY_MATRIX)
	begin	
		if(SEL_MUX_OUTPUT >= 0 and SEL_MUX_OUTPUT < OUTPUT_MUX_SEL_NUMBER) then
			ZERO_FLAG <= ZERO_MATRIX(SEL_MUX_OUTPUT);								   
			CARRY_FLAG <= CARRY_MATRIX(SEL_MUX_OUTPUT);
		else
			ZERO_FLAG <= '0';
			CARRY_FLAG <= '0';
		end if;
	end process;
	
	SECOND_MUX_TAG: MUX_OUTPUT port map(AUXILIAR_MATRIX_OUTPUT, SEL_MUX_OUTPUT, RESULT_OUTPUT);
end architecture ALU_BLACK_BOX_ARCHITECTURE;