entity MICROCONTROLLER_BLACK_BOX is
	


end entity MICROCONTROLLER_BLACK_BOX;